`ifndef AXI4_VIRTUAL_WRITE_SEQ_INCLUDED_
`define AXI4_VIRTUAL_WRITE_SEQ_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: axi4_virtual_write_seq
// Creates and starts the master and slave sequences
//--------------------------------------------------------------------------------------------
class axi4_virtual_write_seq extends uvm_object;
  `uvm_object_utils(axi4_virtual_write_seq)

  //Variable: axi4_master_write_seq_h
  //Instantiation of axi4_master_write_seq handle
  axi4_master_write_seq axi4_master_write_seq_h;

  //Variable: axi4_slave_write_seq_h
  //Instantiation of axi4_slave_write_seq handle
  axi4_slave_write_seq axi4_slave_write_seq_h;

  //-------------------------------------------------------
  // Externally defined Tasks and Functions
  //-------------------------------------------------------
  extern function new(string name = "axi4_virtual_write_seq");
  extern task body();
endclass : axi4_virtual_write_seq

//--------------------------------------------------------------------------------------------
// Construct: new
// Initialises new memory for the object
//
// Parameters:
//  name - axi4_virtual_write_seq
//--------------------------------------------------------------------------------------------
function axi4_virtual_write_seq::new(string name = "axi4_virtual_write_seq");
  super.new(name);
endfunction : new

//--------------------------------------------------------------------------------------------
// Task - body
// Creates and starts the data of master and slave sequences
//--------------------------------------------------------------------------------------------
task axi4_virtual_write_seq::body();
  super.body();
  axi4_master_write_seq_h = axi4_master_write_seq::type_id::create("axi4_master_write_seq_h");
  axi4_slave_write_seq_h = axi4_slave_write_seq::type_id::create("axi4_slave_write_seq_h");
   fork
    forever begin
      axi4_slave_write_seq_h.start(p_sequencer.axi4_slave_seqr_h);
    end
  join_none

  repeat(5) begin
    axi4_master_write_seq_h.start(p_sequencer.axi4_master_seqr_h);
  end
 endtask : body

`endif

