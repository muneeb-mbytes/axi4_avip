`ifndef AXI4_MASTER_NBK_READ_EX_OKAY_RESP_SEQ_INCLUDED_
`define AXI4_MASTER_NBK_READ_EX_OKAY_RESP_SEQ_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: axi4_master_nbk_read_ex_okay_resp_seq
// Extends the axi4_master_nbk_base_seq and randomises the req item
//--------------------------------------------------------------------------------------------
class axi4_master_nbk_read_ex_okay_resp_seq extends axi4_master_nbk_base_seq;
  `uvm_object_utils(axi4_master_nbk_read_ex_okay_resp_seq)

  //-------------------------------------------------------
  // Externally defined Tasks and Functions
  //-------------------------------------------------------
  extern function new(string name = "axi4_master_nbk_read_ex_okay_resp_seq");
  extern task body();
endclass : axi4_master_nbk_read_ex_okay_resp_seq

//--------------------------------------------------------------------------------------------
// Construct: new
// Initializes new memory for the object
//
// Parameters:
//  name - axi4_master_nbk_read_ex_okay_resp_seq
//--------------------------------------------------------------------------------------------
function axi4_master_nbk_read_ex_okay_resp_seq::new(string name = "axi4_master_nbk_read_ex_okay_resp_seq");
  super.new(name);
endfunction : new

//--------------------------------------------------------------------------------------------
// Task: body
// Creates the req of type master_nbk transaction and randomises the req
//--------------------------------------------------------------------------------------------
task axi4_master_nbk_read_ex_okay_resp_seq::body();
  super.body();
  req.transfer_type=NON_BLOCKING_READ;
//  req = axi4_master_nbk_tx::type_id::create("req");
  //req.axi4_master_nbk_agent_cfg_h = p_sequencer.axi4_master_nbk_agent_cfg_h;
  
  start_item(req);
  if(!req.randomize() with {req.arsize == READ_4_BYTES;
                            req.tx_type == READ;
                            req.arburst == READ_INCR;
                            req.transfer_type == NON_BLOCKING_READ;}) begin

    `uvm_fatal("axi4","Rand failed");
  end
  req.print();
  finish_item(req);
endtask : body

`endif

